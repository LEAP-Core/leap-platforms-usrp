Bit#(32) samples[1024] = {
32'hdeaddead,
32'hcafecafe,
32'h02f102f1,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h020f020f,
32'h001afa11,
32'hfc7bff65,
32'hff6e0664,
32'h0000041e,
32'hff6e0664,
32'hfc7bff65,
32'h001afa11,
32'h020f020f,
32'hfa11001a,
32'hff65fc7b,
32'h0664ff6e,
32'h041e0000,
32'h0664ff6e,
32'hff65fc7b,
32'hfa11001a,
32'h0000f900,
32'hfba0008c,
32'hfb41041b,
32'hfad7fbe1,
32'hfd97ffdf,
32'h0351035c,
32'h00eafa4b,
32'h00bdfa89,
32'h06c2fe6d,
32'h00f9fd77,
32'hfc5bfd4b,
32'hff5d031d,
32'hfbdc03ae,
32'hfd13fa1e,
32'hfe3dfd6f,
32'hfb9701a6,
32'h02cc02cc,
32'h002e0557,
32'hf8cdfefd,
32'h00aa02a0,
32'h029e0118,
32'h021ff9de,
32'h0526000b,
32'hffd10263,
32'h0128045e,
32'h04c1fe48,
32'h0278fad7,
32'h03ed02ad,
32'hfec000f1,
32'hfc4a0456,
32'h04fa01c7,
32'h0563ffc5,
32'h000006ff,
32'hfa9bffc5,
32'hfb0401c7,
32'h03b50456,
32'h013f00f1,
32'hfc1102ad,
32'hfd86fad7,
32'hfb3efe48,
32'hfed6045e,
32'h002e0263,
32'hfad8000b,
32'hfde0f9de,
32'hfd600118,
32'hff5402a0,
32'h0732fefd,
32'hffd00557,
32'hfd3302cc,
32'h046701a6,
32'h01c2fd6f,
32'h02ebfa1e,
32'h042303ae,
32'h00a1031d,
32'h03a3fd4b,
32'hff05fd77,
32'hf93dfe6d,
32'hff41fa89,
32'hff14fa4b,
32'hfcae035c,
32'h0267ffdf,
32'h0528fbe1,
32'h04bd041b,
32'h045f008c,
32'h0000f900,
32'hfba0008c,
32'hfb41041b,
32'hfad7fbe1,
32'hfd97ffdf,
32'h0351035c,
32'h00eafa4b,
32'h00bdfa89,
32'h06c2fe6d,
32'h00f9fd77,
32'hfc5bfd4b,
32'hff5d031d,
32'hfbdc03ae,
32'hfd13fa1e,
32'hfe3dfd6f,
32'hfb9701a6,
32'h02cc02cc,
32'h002e0557,
32'hf8cdfefd,
32'h00aa02a0,
32'h029e0118,
32'h021ff9de,
32'h0526000b,
32'hffd10263,
32'h0128045e,
32'h04c1fe48,
32'h0278fad7,
32'h03ed02ad,
32'hfec000f1,
32'hfc4a0456,
32'h04fa01c7,
32'h0563ffc5,
32'h000006ff,
32'hfa9bffc5,
32'hfb0401c7,
32'h03b50456,
32'h013f00f1,
32'hfc1102ad,
32'hfd86fad7,
32'hfb3efe48,
32'hfed6045e,
32'h002e0263,
32'hfad8000b,
32'hfde0f9de,
32'hfd600118,
32'hff5402a0,
32'h0732fefd,
32'hffd00557,
32'hfd3302cc,
32'h046701a6,
32'h01c2fd6f,
32'h02ebfa1e,
32'h042303ae,
32'h00a1031d,
32'h03a3fd4b,
32'hff05fd77,
32'hf93dfe6d,
32'hff41fa89,
32'hff14fa4b,
32'hfcae035c,
32'h0267ffdf,
32'h0528fbe1,
32'h04bd041b,
32'h045f008c,
32'h0000f900,
32'hfba0008c,
32'hfb41041b,
32'hfad7fbe1,
32'hfd97ffdf,
32'h0351035c,
32'h00eafa4b,
32'h00bdfa89,
32'h06c2fe6d,
32'h00f9fd77,
32'hfc5bfd4b,
32'hff5d031d,
32'hfbdc03ae,
32'hfd13fa1e,
32'hfe3dfd6f,
32'hfb9701a6,
32'h02cc02cc,
32'h002e0557,
32'hf8cdfefd,
32'h00aa02a0,
32'h029e0118,
32'h021ff9de,
32'h0526000b,
32'hffd10263,
32'h0128045e,
32'h04c1fe48,
32'h0278fad7,
32'h03ed02ad,
32'hfec000f1,
32'hfc4a0456,
32'h04fa01c7,
32'h0563ffc5,
32'hffff0166,
32'hfe9705c4,
32'hfa990210,
32'hffa9029f,
32'h03760154,
32'h05b8fad3,
32'h0404fddb,
32'hff4d00d1,
32'h028e045d,
32'h013ffd62,
32'h010bfb8b,
32'h05f804a3,
32'hfd0001c9,
32'hfd6204f9,
32'h08cf01bf,
32'h03e1fe91,
32'hfffd0598,
32'hfc1efe91,
32'hf73001bd,
32'h029c04f9,
32'h02fd01c9,
32'hfa0504a1,
32'hfef3fb8a,
32'hfec1fd63,
32'hfd70045d,
32'h00b100d1,
32'hfbf9fddb,
32'hfa47fad0,
32'hfc890154,
32'h0055029f,
32'h05650211,
32'h016605c4,
32'h00000165,
32'h03a902c7,
32'h028dfb6f,
32'h0361f75f,
32'h0150056e,
32'hffc702b6,
32'h03b3fce4,
32'hfdf9015d,
32'hfaa4fe6c,
32'h0136f91b,
32'hff6ffc2e,
32'hfd6100db,
32'h022cfd0d,
32'h0384fdfd,
32'h037f0311,
32'h038d0031,
32'h0000fd33,
32'hfc710031,
32'hfc7f0310,
32'hfc7cfdfd,
32'hfdd2fd0e,
32'h029d00db,
32'h0090fc2f,
32'hfec9f91a,
32'h055bfe6e,
32'h0205015f,
32'hfc4cfce4,
32'h003702b6,
32'hfeae056d,
32'hfca0f75e,
32'hfd72fb6f,
32'hfc5502c7,
32'hffff0166,
32'hfe9705c4,
32'hfa990210,
32'hffa9029f,
32'h03760154,
32'h05b8fad3,
32'h0404fddb,
32'hff4d00d1,
32'h028e045d,
32'h013ffd62,
32'h010bfb8b,
32'h05f804a3,
32'hfd0001c9,
32'hfd6204f9,
32'h08cf01bf,
32'h03e1fe91,
32'hfcc200c8,
32'hfb52010a,
32'h0117008b,
32'hfe80ff3d,
32'hfcd40277,
32'hfbf4026f,
32'hfa11fee8,
32'hfe60feab,
32'h0005fd90,
32'hfb3ffe0c,
32'hfcf4ffbc,
32'h047200d4,
32'h00c60320,
32'hfbf70122,
32'hffc800b1,
32'hfeec01cf,
32'hfe73fe39,
32'h00d0fb7d,
32'h011afc79,
32'h01a30312,
32'h00620267,
32'hff19f9fc,
32'hff6dfea4,
32'h018f04d6,
32'h0109014e,
32'hfec2fd10,
32'hff72fc5b,
32'hfe030001,
32'h01b700bf,
32'h0449ffe4,
32'hfdcc018e,
32'hffa100d4,
32'h01cbfed1,
32'hfec5fe24,
32'h0320fe4c,
32'h043afec0,
32'hfd0c0206,
32'hfe05047b,
32'h03d90332,
32'hfe0a0257,
32'hfe72ff53,
32'h0634ffcd,
32'h00bb0278,
32'h0231fead,
32'h0503fd66,
32'hfb19fec0,
32'hfd91004a,
32'h04e90203,
32'h02a4026d,
32'hffa303db,
32'hfe6efe62,
32'hffe1fa24,
32'h00eafcc3,
32'hff6efbc1,
32'h0030ffb8,
32'h03a70401,
32'h023d00a8,
32'hfe32ff1e,
32'hfe93fef9,
32'h0096010e,
32'h03f201e0,
32'h025efe5d,
32'hffc8ffc6,
32'h022c024d,
32'hfcc200c8,
32'hfb52010a,
32'h0117008b,
32'hfe80ff3d,
32'hfcd40277,
32'hfbf4026f,
32'hfa11fee8,
32'hfe60feab,
32'h0005fd90,
32'hfb3ffe0c,
32'hfcf4ffbc,
32'h047200d4,
32'h00c60320,
32'hfbf70122,
32'hffc800b1,
32'hfeec01cf,
32'h0030040b,
32'h02d4fead,
32'hff1ffece,
32'hfe5cfd0d,
32'hff2b0075,
32'hfe7f042a,
32'hfda8ffa4,
32'h033501bd,
32'h0464000c,
32'hfb01fd04,
32'hfeec0454,
32'h04970395,
32'hff760012,
32'h01fc0259,
32'h02fc004d,
32'hfc56fc69,
32'hfcf0fb01,
32'h02050118,
32'h01e604d4,
32'h006d002c,
32'hff92026d,
32'hfe620106,
32'hffd3fd18,
32'h011b024e,
32'h035400b1,
32'h02870066,
32'h002d01e5,
32'h0443fd8e,
32'h00f10213,
32'hfe33038c,
32'h011901a6,
32'hfd2e02d5,
32'h0097fd43,
32'h016bfcfe,
32'hfe90fd78,
32'h043bfb06,
32'hfdf0fdf3,
32'hf9e8fd0e,
32'h01a5feab,
32'h013a030c,
32'hff68029d,
32'hff740098,
32'hff00fe2d,
32'hffd10022,
32'hffb9feb0,
32'hfdf9fd71,
32'hfdcb046b,
32'h02d10338,
32'h03520086,
32'hffa70431,
32'hfed40282,
32'hfc3fff05,
32'hfc7dfd67,
32'hfee8fba7,
32'hfd46fc64,
32'hfe8fffbb,
32'h0142ff9c,
32'hfc74fe57,
32'hfd57fef7,
32'h0644fd40,
32'h02240114,
32'hfe6601c3,
32'h02effad2,
32'hffac008d,
32'h0030040b,
32'h02d4fead,
32'hff1ffece,
32'hfe5cfd0d,
32'hff2b0075,
32'hfe7f042a,
32'hfda8ffa4,
32'h033501bd,
32'h0464000c,
32'hfb01fd04,
32'hfeec0454,
32'h04970395,
32'hff760012,
32'h01fc0259,
32'h02fc004d,
32'hfc56fc69,
32'hfe1eff19,
32'h00b1fe97,
32'h047b0037,
32'hff20045b,
32'hfddf0467,
32'h00bffd91,
32'hfcf9fa57,
32'h0125fe01,
32'h023f0236,
32'hff0b022f,
32'h00cf0090,
32'h001f0092,
32'h026a006f,
32'h0206ff2e,
32'hfe63fead,
32'hfde2ff48,
32'hff4cff72,
32'h00c7fd8e,
32'hfc63fb70,
32'hfe0a005b,
32'h005802fd,
32'hfc7cff5a,
32'hfedf05c9,
32'hfc6e0607,
32'hfc1af959,
32'h0170f86f,
32'h000dfef3,
32'h01590482,
32'h022b056e,
32'h0068ffa9,
32'hfe35fdb1,
32'h0000fe94,
32'h06080097,
32'hfeb50244,
32'hfb48005f,
32'h012dfd79,
32'hfbd2fde2,
32'hfb5c01e9,
32'h0120ff20,
32'hffd9fd91,
32'hff47008b,
32'h0198fe51,
32'h02ea020a,
32'h0392013a,
32'h049cfb78,
32'h02dd025c,
32'h0140044e,
32'h038500d6,
32'h012d0133,
32'hfd6d007d,
32'h02a200c3,
32'h0427fe86,
32'hfd8efd12,
32'h001efead,
32'h022bff0d,
32'hfd16fee2,
32'hff220037,
32'hfff903bc,
32'hff58014b,
32'hffb3ff99,
32'hfd710378,
32'h00e70014,
32'h016bfd80,
32'hfe34ffc4,
32'hfe1eff19,
32'h00b1fe97,
32'h047b0037,
32'hff20045b,
32'hfddf0467,
32'h00bffd91,
32'hfcf9fa57,
32'h0125fe01,
32'h023f0236,
32'hff0b022f,
32'h00cf0090,
32'h001f0092,
32'h026a006f,
32'h0206ff2e,
32'hfe63fead,
32'hfde2ff48,
32'h046a01af,
32'h0166011c,
32'h02a2ff9f,
32'hff46fd47,
32'hfd1effcf,
32'hffb3ff4e,
32'h006a01a3,
32'hfffd01e9,
32'hfd38fd4c,
32'h012cfdf3,
32'h00fa00d6,
32'hfdd901d2,
32'h0149fe60,
32'hffeaffa5,
32'h00ed04e5,
32'h0133041e,
32'h002c0357,
32'h01f8ff68,
32'hff9ffe40,
32'h00350085,
32'hff06fc57,
32'hffb1fe03,
32'h01adff52,
32'hff35fedd,
32'h042a0481,
32'h00ce005d,
32'hfbc0fd1f,
32'h032e03bb,
32'h018002a6,
32'hfbe5fe49,
32'hfc4bfe76,
32'hffc8ff7c,
32'h02ab003d,
32'h0127fe54,
32'hfec7fe10,
32'hfd0c02d9,
32'h01020201,
32'h026afd80,
32'hfe27feba,
32'h0031ff5d,
32'h016cff27,
32'h013000f4,
32'h057a0169,
32'h04d30064,
32'hfce6ff1a,
32'hfdd2ff82,
32'h0481ff02,
32'h0263fe46,
32'h0289fde0,
32'hff38fd1d,
32'hf9f30042,
32'h0026ffe9,
32'hff29fdfc,
32'hfbc9018a,
32'hfd03038d,
32'hfd31021d,
32'hff76fb88,
32'hfe71f9a6,
32'h00b2000a,
32'hfec4011d,
32'hfbc00035,
32'h0201ffca,
32'hff3e0299,
32'h001b05b8,
32'h046a01af,
32'h0166011c,
32'h02a2ff9f,
32'hff46fd47,
32'hfd1effcf,
32'hffb3ff4e,
32'h006a01a3,
32'hfffd01e9,
32'hfd38fd4c,
32'h012cfdf3,
32'h00fa00d6,
32'hfdd901d2,
32'h0149fe60,
32'hffeaffa5,
32'h00ed04e5,
32'h0133041e,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h0000000f};
