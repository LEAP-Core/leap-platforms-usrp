typedef 2048 NumSamples;
typedef 1363 PacketLength;

Bit#(32) samples[2048] = {
32'hdeaddead,
32'hcafecafe,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'hf6000000,
32'h00c9f9c0,
32'h05def939,
32'hfa1ef8a1,
32'hffd1fc8f,
32'h04cd04bd,
32'hf7d9014f,
32'hf832010f,
32'hfdc109a8,
32'hfc620165,
32'hfc23facc,
32'h0473ff18,
32'h0543fa16,
32'hf799fbd3,
32'hfc56fd7c,
32'h025cf9b4,
32'h04000400,
32'h07a10043,
32'hfe8ff5b7,
32'h03c100f4,
32'h019103be,
32'hf73e0308,
32'h0010075c,
32'h0369ffbd,
32'h063e01a8,
32'hfd8c06cb,
32'hf8a10388,
32'h03d4059d,
32'h0159fe37,
32'h0632fab3,
32'h028b071d,
32'hffac07b3,
32'h0a000000,
32'hffacf84c,
32'h028bf8e2,
32'h0632054c,
32'h015901c8,
32'h03d4fa62,
32'hf8a1fc77,
32'hfd8cf934,
32'h063efe57,
32'h03690042,
32'h0010f8a3,
32'hf73efcf7,
32'h0191fc41,
32'h03c1ff0b,
32'hfe8f0a48,
32'h07a1ffbc,
32'h0400fc00,
32'h025c064b,
32'hfc560283,
32'hf799042c,
32'h054305e9,
32'h047300e7,
32'hfc230533,
32'hfc62fe9a,
32'hfdc1f657,
32'hf832fef0,
32'hf7d9feb0,
32'h04cdfb42,
32'hffd10370,
32'hfa1e075e,
32'h05de06c6,
32'h00c9063f,
32'hf6000000,
32'h00c9f9c0,
32'h05def939,
32'hfa1ef8a1,
32'hffd1fc8f,
32'h04cd04bd,
32'hf7d9014f,
32'hf832010f,
32'hfdc109a8,
32'hfc620165,
32'hfc23facc,
32'h0473ff18,
32'h0543fa16,
32'hf799fbd3,
32'hfc56fd7c,
32'h025cf9b4,
32'h04000400,
32'h07a10043,
32'hfe8ff5b7,
32'h03c100f4,
32'h019103be,
32'hf73e0308,
32'h0010075c,
32'h0369ffbd,
32'h063e01a8,
32'hfd8c06cb,
32'hf8a10388,
32'h03d4059d,
32'h0159fe37,
32'h0632fab3,
32'h028b071d,
32'hffac07b3,
32'h0a000000,
32'hffacf84c,
32'h028bf8e2,
32'h0632054c,
32'h015901c8,
32'h03d4fa62,
32'hf8a1fc77,
32'hfd8cf934,
32'h063efe57,
32'h03690042,
32'h0010f8a3,
32'hf73efcf7,
32'h0191fc41,
32'h03c1ff0b,
32'hfe8f0a48,
32'h07a1ffbc,
32'h0400fc00,
32'h025c064b,
32'hfc560283,
32'hf799042c,
32'h054305e9,
32'h047300e7,
32'hfc230533,
32'hfc62fe9a,
32'hfdc1f657,
32'hf832fef0,
32'hf7d9feb0,
32'h04cdfb42,
32'hffd10370,
32'hfa1e075e,
32'h05de06c6,
32'h00c9063f,
32'hf6000000,
32'h00c9f9c0,
32'h05def939,
32'hfa1ef8a1,
32'hffd1fc8f,
32'h04cd04bd,
32'hf7d9014f,
32'hf832010f,
32'hfdc109a8,
32'hfc620165,
32'hfc23facc,
32'h0473ff18,
32'h0543fa16,
32'hf799fbd3,
32'hfc56fd7c,
32'h025cf9b4,
32'h04000400,
32'h07a10043,
32'hfe8ff5b7,
32'h03c100f4,
32'h019103be,
32'hf73e0308,
32'h0010075c,
32'h0369ffbd,
32'h063e01a8,
32'hfd8c06cb,
32'hf8a10388,
32'h03d4059d,
32'h0159fe37,
32'h0632fab3,
32'h028b071d,
32'hffac07b3,
32'h0200ffff,
32'h083dfdfd,
32'h02f3f849,
32'h03c0ff84,
32'h01e604f2,
32'hf89c082c,
32'hfcf105bd,
32'h012cff01,
32'h063d03a7,
32'hfc4301c8,
32'hf9a2017e,
32'h06a00888,
32'h028dfbb7,
32'h071cfc43,
32'h02800c96,
32'hfdf5058b,
32'h07fefffd,
32'hfdf4fa75,
32'h027df36a,
32'h071c03bb,
32'h028d0446,
32'h069df775,
32'hf9a1fe81,
32'hfc45fe39,
32'h063dfc57,
32'h012c00fd,
32'hfcf0fa40,
32'hf898f7d4,
32'h01e6fb0e,
32'h03c0007a,
32'h02f407b6,
32'h083e0200,
32'h01ff0000,
32'h03f8053c,
32'hf97b03a5,
32'hf3ad04d5,
32'h07c201e1,
32'h03e0ffaf,
32'hfb900549,
32'h01f3fd1b,
32'hfdc0f858,
32'hf62701bc,
32'hfa8cff32,
32'h013afc42,
32'hfbca031b,
32'hfd210506,
32'h046204ff,
32'h00470514,
32'hfc000000,
32'h0047faeb,
32'h0461faff,
32'hfd21fafb,
32'hfbcbfce4,
32'h013903bc,
32'hfa8d00ce,
32'hf626fe44,
32'hfdc307a7,
32'h01f602e4,
32'hfb8ffab6,
32'h03e00050,
32'h07c1fe1e,
32'hf3acfb2e,
32'hf97bfc5b,
32'h03f8fac3,
32'h0200ffff,
32'h083dfdfd,
32'h02f3f849,
32'h03c0ff84,
32'h01e604f2,
32'hf89c082c,
32'hfcf105bd,
32'h012cff01,
32'h063d03a7,
32'hfc4301c8,
32'hf9a2017e,
32'h06a00888,
32'h028dfbb7,
32'h071cfc43,
32'h02800c96,
32'hfdf5058b,
32'h011efb5f,
32'h017df951,
32'h00c70190,
32'hfeeafddc,
32'h0386fb79,
32'h037bfa39,
32'hfe70f786,
32'hfe19fdae,
32'hfc850008,
32'hfd36f936,
32'hffa0fba6,
32'h0130065b,
32'h0477011c,
32'h019ffa3d,
32'h00feffb0,
32'h0296fe76,
32'hfd76fdc9,
32'hf98f012a,
32'hfaf60194,
32'h04630258,
32'h0370008d,
32'hf768feb6,
32'hfe0fff2e,
32'h06e9023b,
32'h01de017b,
32'hfbcffe3b,
32'hfaccff36,
32'h0002fd2a,
32'h01120274,
32'hffd90620,
32'h0239fcdb,
32'h0130ff79,
32'hfe500290,
32'hfd59fe3e,
32'hfd920478,
32'hfe38060a,
32'h02e5fbc8,
32'h0668fd2c,
32'h04910580,
32'h0358fd34,
32'hff0afdc8,
32'hffb808dd,
32'h0387010c,
32'hfe1c0322,
32'hfc490729,
32'hfe38f900,
32'h006bfc87,
32'h02e10705,
32'h037803c6,
32'h0583ff7c,
32'hfdb1fdc2,
32'hf7a2ffd5,
32'hfb61014f,
32'hf9f0ff30,
32'hff9a0046,
32'h05b90539,
32'h00f10333,
32'hfebefd6d,
32'hfe89fdf7,
32'h018300d7,
32'h02af05a4,
32'hfdaa0362,
32'hffaeffb0,
32'h034a031b,
32'h011efb5f,
32'h017df951,
32'h00c70190,
32'hfeeafddc,
32'h0386fb79,
32'h037bfa39,
32'hfe70f786,
32'hfe19fdae,
32'hfc850008,
32'hfd36f936,
32'hffa0fba6,
32'h0130065b,
32'h0477011c,
32'h019ffa3d,
32'h00feffb0,
32'h0296fe76,
32'h05c70046,
32'hfe1c040b,
32'hfe4bfebf,
32'hfbcafda9,
32'h00a8fed1,
32'h05f4fdda,
32'hff7dfca7,
32'h027d0495,
32'h00120646,
32'hfbbdf8de,
32'h062ffe77,
32'h051f0690,
32'h001bff3b,
32'h035c02d7,
32'h006f0444,
32'hfae0fac4,
32'hf8defba1,
32'h019102e4,
32'h06e602b7,
32'h003f009c,
32'h0378ff64,
32'h0177fdb1,
32'hfbdaffc1,
32'h034b0195,
32'h00fe04c2,
32'h0093039d,
32'h02b60041,
32'hfc820618,
32'h02f80159,
32'h0512fd6e,
32'h025c0192,
32'h040dfbf9,
32'hfc1700d8,
32'hfbb40208,
32'hfc63fdf3,
32'hf8e4060c,
32'hfd13fd0f,
32'hfbcbf74c,
32'hfe19025a,
32'h045b01c2,
32'h03bdff28,
32'h00daff38,
32'hfd66fe93,
32'h0032ffbd,
32'hfe21ff9b,
32'hfc59fd1b,
32'h0651fcda,
32'h049a0407,
32'h00c004bf,
32'h05fdff82,
32'h0396fe54,
32'hfe9afaa4,
32'hfc4afafc,
32'hf9cafe70,
32'hfad8fc1b,
32'hff9efdf1,
32'hff7201cd,
32'hfda2faef,
32'hfe86fc34,
32'hfc1308f4,
32'h018b030f,
32'h0285fdb7,
32'hf89a0432,
32'h00caff89,
32'h05c70046,
32'hfe1c040b,
32'hfe4bfebf,
32'hfbcafda9,
32'h00a8fed1,
32'h05f4fdda,
32'hff7dfca7,
32'h027d0495,
32'h00120646,
32'hfbbdf8de,
32'h062ffe77,
32'h051f0690,
32'h001bff3b,
32'h035c02d7,
32'h006f0444,
32'hfae0fac4,
32'hfeb7fd50,
32'hfdfd00fd,
32'h004f0668,
32'h063afec0,
32'h064bfcf6,
32'hfc860112,
32'hf7eafbae,
32'hfd2701a3,
32'h03290336,
32'h0320fea3,
32'h00ce0129,
32'h00d1002d,
32'h009f0374,
32'hfed502e5,
32'hfe1dfdb2,
32'hfefafcfa,
32'hff36ff00,
32'hfc82011d,
32'hf97cfad7,
32'h0083fd34,
32'h0446007e,
32'hff14fafb,
32'h0844fe64,
32'h089dfae7,
32'hf67ffa6f,
32'hf531020f,
32'hfe810014,
32'h067201ee,
32'h07c20319,
32'hff840096,
32'hfcb5fd71,
32'hfdf80000,
32'h00d9089f,
32'h033dfe28,
32'h0088f943,
32'hfc6501af,
32'hfcfafa08,
32'h02bbf95f,
32'hfec1019c,
32'hfc86ffc9,
32'h00c7fef8,
32'hfd990247,
32'h02eb042a,
32'h01c1051a,
32'hf9880697,
32'h035f0418,
32'h062701ca,
32'h01330508,
32'h01b701af,
32'h00b3fc53,
32'h011803c3,
32'hfde405f0,
32'hfbd1fc82,
32'hfe1c002b,
32'hfea6031a,
32'hfe68fbd7,
32'h004ffec3,
32'h0557fff7,
32'h01daff10,
32'hff6dff93,
32'h04f5fc59,
32'h001e014b,
32'hfc6e0207,
32'hffabfd6f,
32'hfeb7fd50,
32'hfdfd00fd,
32'h004f0668,
32'h063afec0,
32'h064bfcf6,
32'hfc860112,
32'hf7eafbae,
32'hfd2701a3,
32'h03290336,
32'h0320fea3,
32'h00ce0129,
32'h00d1002d,
32'h009f0374,
32'hfed502e5,
32'hfe1dfdb2,
32'hfefafcfa,
32'h0268064f,
32'h01960200,
32'hff7603c3,
32'hfc1dfef7,
32'hffbafbe3,
32'hff02ff92,
32'h02570098,
32'h02bbfffd,
32'hfc24fc07,
32'hfd1301ad,
32'h01320166,
32'h029afced,
32'hfdae01d7,
32'hff7fffe1,
32'h06ff0153,
32'h05e301b8,
32'h04c6003f,
32'hff2802d1,
32'hfd81ff76,
32'h00bf004c,
32'hfac6fe9c,
32'hfd29ff90,
32'hff080266,
32'hfe61fedf,
32'h067005f3,
32'h00860127,
32'hfbe4f9ee,
32'h0555048b,
32'h03ca0226,
32'hfd8efa23,
32'hfdcefab5,
32'hff44ffb1,
32'h005803d0,
32'hfd9d01a6,
32'hfd3cfe41,
32'h0412fbc8,
32'h02de0172,
32'hfc6e0374,
32'hfe2ffd5d,
32'hff180047,
32'hfecb0209,
32'h015d01b3,
32'h020507d4,
32'h008f06e5,
32'hfeb8fb92,
32'hff4dfce3,
32'hfe960670,
32'hfd890369,
32'hfcf803a0,
32'hfbe1fee3,
32'h005ff75b,
32'hffe00037,
32'hfd20fece,
32'h0234f9fb,
32'h0513fbbc,
32'h0305fbfe,
32'hf99fff3c,
32'hf6eefdc6,
32'h000f00ff,
32'h0198fe3d,
32'h004df9ef,
32'hffb302dd,
32'h03b7feec,
32'h082c0027,
32'h0268064f,
32'h01960200,
32'hff7603c3,
32'hfc1dfef7,
32'hffbafbe3,
32'hff02ff92,
32'h02570098,
32'h02bbfffd,
32'hfc24fc07,
32'hfd1301ad,
32'h01320166,
32'h029afced,
32'hfdae01d7,
32'hff7fffe1,
32'h06ff0153,
32'h05e301b8,
32'h0380010f,
32'h0009fcb2,
32'hfa37026b,
32'hfd50028e,
32'hfeabfc36,
32'hfa98ffd6,
32'hfcee0152,
32'h048f0001,
32'h071401a2,
32'hff6dff84,
32'hf9b2fffa,
32'hfc3d05e4,
32'hfa34058a,
32'hfd12fe1f,
32'h0252fb6e,
32'hfccffcc5,
32'h0086fc08,
32'h02c2fd8a,
32'hfd5000db,
32'h00830184,
32'hfc7a0295,
32'hf97a06c4,
32'hfdb90694,
32'hfe64015a,
32'h01d800f5,
32'h021200d2,
32'h003000da,
32'hfcdc053f,
32'hfb59021a,
32'hff59fa28,
32'h0055f8ef,
32'h04cefb2e,
32'h034ffbbf,
32'h0727fd10,
32'h11490044,
32'h004eff16,
32'hfaf3fddf,
32'h055dfe6a,
32'hfffcfda5,
32'h01560353,
32'hfdab02bd,
32'hf971fa94,
32'h01a20129,
32'h01660547,
32'h0083fc61,
32'hfdf3ffa8,
32'hfadf059a,
32'h01b0fcba,
32'h0727fca6,
32'h0416063c,
32'hfefc016a,
32'h034fff0f,
32'h04a60615,
32'h024701b3,
32'h06d4fda6,
32'h02f8fece,
32'h00a6f9aa,
32'h0005fb7c,
32'hf76d018c,
32'hfd2afe5f,
32'h04efffba,
32'hfe680367,
32'hfac0ff53,
32'hfed300cd,
32'h0380010f,
32'h0009fcb2,
32'hfa37026b,
32'hfd50028e,
32'hfeabfc36,
32'hfa98ffd6,
32'hfcee0152,
32'h048f0001,
32'h071401a2,
32'hff6dff84,
32'hf9b2fffa,
32'hfc3d05e4,
32'hfa34058a,
32'hfd12fe1f,
32'h0252fb6e,
32'hfccffcc5,
32'hfc210320,
32'h01a00431,
32'h001900b5,
32'hfd52f730,
32'hfedefa15,
32'hfbd2fd7a,
32'hfafa00be,
32'h02e50074,
32'h051ffc37,
32'hfe56032c,
32'h0156012a,
32'h0821fd76,
32'h038c05c2,
32'h00410717,
32'h024c0186,
32'h060afdb0,
32'h0695fb46,
32'h014ff9c3,
32'h00c601db,
32'hfb290166,
32'hf70df877,
32'h02db0281,
32'h047100cf,
32'h005afc0d,
32'h03bf05fe,
32'hff8bffd9,
32'hfec0feaa,
32'h025affa5,
32'hff86f9b5,
32'h0028003d,
32'hfd1c01cd,
32'hf6ecffaa,
32'hfe40ffe0,
32'h03db0395,
32'h02d80734,
32'h0663fe7d,
32'h03e40023,
32'hff80061a,
32'hfaf4009f,
32'hf83b00c8,
32'h04cf0097,
32'h04d3fd65,
32'hf7c4014c,
32'hfa8002ef,
32'h00eaff2a,
32'h063d036d,
32'h01fc031b,
32'hf897f913,
32'hfe87fe38,
32'hfeb702fb,
32'hfceafeba,
32'h025b023b,
32'hfd4d0231,
32'hfcc0fd16,
32'h02dffd31,
32'h00cd0461,
32'hfa1205f2,
32'hf62bfe12,
32'hfe01fbdf,
32'h04eefeac,
32'h0123043b,
32'h0384000a,
32'h0758f7b1,
32'hff80fedc,
32'hfc210320,
32'h01a00431,
32'h001900b5,
32'hfd52f730,
32'hfedefa15,
32'hfbd2fd7a,
32'hfafa00be,
32'h02e50074,
32'h051ffc37,
32'hfe56032c,
32'h0156012a,
32'h0821fd76,
32'h038c05c2,
32'h00410717,
32'h024c0186,
32'h060afdb0,
32'h06a00106,
32'h03ba0618,
32'hf97001ab,
32'h0065fc34,
32'hfebd0116,
32'hfdf6038c,
32'h034700bd,
32'hfb89fdfc,
32'hffba02f4,
32'h00eb00c3,
32'hff67fa21,
32'h048fffd5,
32'h023400ca,
32'h076d03e9,
32'h025f082b,
32'hfed5ff1a,
32'h055dfb47,
32'hfc29feba,
32'hff8a021f,
32'h0235ffbd,
32'hfd07fab3,
32'h0323fbc4,
32'hfe18fd98,
32'hfc03017a,
32'hfe4cff42,
32'hfc80fda2,
32'h009ffd99,
32'hfd7ef3b7,
32'hffe5fb96,
32'h09540453,
32'h04adfca7,
32'hffe00054,
32'h02900308,
32'hfd1c01dc,
32'hf768ff97,
32'hfce2fa8f,
32'hfe5eff40,
32'hff0f02d5,
32'h02e3030f,
32'h0226feb1,
32'h0315fb5b,
32'h0173029f,
32'h001cff35,
32'hff86fa8d,
32'hfdd8010f,
32'h009d0206,
32'hff9f0254,
32'h02ba032b,
32'h038ffe67,
32'hff26fddb,
32'h045601a3,
32'hff65ff83,
32'hf73c0138,
32'hfa860840,
32'hfe0a0444,
32'hff750288,
32'hfc4406ae,
32'hfeb6fecd,
32'h0261fa4a,
32'hfebb02a6,
32'hfdae014f,
32'hffb7f9f5,
32'h0148ffec,
32'h00b202f1,
32'h06a00106,
32'h03ba0618,
32'hf97001ab,
32'h0065fc34,
32'hfebd0116,
32'hfdf6038c,
32'h034700bd,
32'hfb89fdfc,
32'hffba02f4,
32'h00eb00c3,
32'hff67fa21,
32'h048fffd5,
32'h023400ca,
32'h076d03e9,
32'h025f082b,
32'hfed5ff1a,
32'hfc900358,
32'hfca6f977,
32'hfe1efbfe,
32'hfbf10c2b,
32'hfc3302a6,
32'hffe2fb04,
32'h015b0021,
32'h0506fe0a,
32'h064cfd20,
32'hfe3f029f,
32'hfb6c0782,
32'hff7fffb0,
32'hfd80fbbf,
32'hfb30fe3d,
32'hfdc4fc76,
32'hfcc0016b,
32'hfe36fc60,
32'h0540f9b1,
32'h035b0340,
32'hffec0265,
32'h00ac0279,
32'hfd6bfd69,
32'hfea4fd43,
32'h0030085b,
32'hff88040d,
32'h068a014c,
32'h04a7003c,
32'hf813fd4d,
32'hf8c000d8,
32'h0116ff4e,
32'h024a002b,
32'h0104ff6a,
32'h01d00217,
32'h05720600,
32'h0403fb28,
32'hfd49fe4c,
32'hff4705cf,
32'hfef1fbb0,
32'hfc09f7b0,
32'h02ddfe3d,
32'h019201ae,
32'hfdb4f94a,
32'h00cbfa61,
32'hff940757,
32'hfd3200b2,
32'hfbbdfcaa,
32'h010e04cf,
32'h00bf00cf,
32'hf9280231,
32'h01740616,
32'h00f2fd44,
32'hfcabfdbf,
32'h0899ffce,
32'h062cfb18,
32'h026f0368,
32'h06070773,
32'h0157fee1,
32'h00fbfac6,
32'hfd6efb33,
32'hfa5c0198,
32'h024c0636,
32'h04c402d5,
32'h02a8fd0f,
32'h008bfe38,
32'hfc900358,
32'hfca6f977,
32'hfe1efbfe,
32'hfbf10c2b,
32'hfc3302a6,
32'hffe2fb04,
32'h015b0021,
32'h0506fe0a,
32'h064cfd20,
32'hfe3f029f,
32'hfb6c0782,
32'hff7fffb0,
32'hfd80fbbf,
32'hfb30fe3d,
32'hfdc4fc76,
32'hfcc0016b,
32'h00b905df,
32'hffa200df,
32'hf85dffcf,
32'hfed30752,
32'h000dfcec,
32'hfff7fcf6,
32'h03a90286,
32'h0296fe8b,
32'h011003dc,
32'h03780419,
32'h038e019a,
32'hfba30046,
32'hfc10fec0,
32'h015a027b,
32'h013fff87,
32'h026a0477,
32'hff07028f,
32'h015bf6dd,
32'h02f8007e,
32'hfabaffad,
32'hfb03f9e0,
32'hf807fee7,
32'hf888fd8e,
32'h059904d7,
32'h049a05d6,
32'hfe65005c,
32'h0072016b,
32'h00bb00b6,
32'h00ad0500,
32'h006e01c2,
32'hfcdf012f,
32'h01020467,
32'h0806fbde,
32'h051e0140,
32'h046b03e3,
32'hffdbfb70,
32'hfc820055,
32'h0669011b,
32'h010bfe34,
32'hf891014f,
32'hfbf0ff43,
32'hfcc1fe86,
32'h01540185,
32'h00f1f7a5,
32'h0089f214,
32'h02140069,
32'hfe4efe58,
32'h03c8f6e6,
32'h0237fed0,
32'hfc17fb38,
32'h00ccfc17,
32'hfe8f02a3,
32'hfc6cff7f,
32'h03110249,
32'h061b019f,
32'h00630134,
32'hfe2602a8,
32'h0301fca2,
32'hff1c0329,
32'hfb37048c,
32'h0276f9cb,
32'h0752013e,
32'hfdba0407,
32'hf6a6ff0f,
32'h00b905df,
32'hffa200df,
32'hf85dffcf,
32'hfed30752,
32'h000dfcec,
32'hfff7fcf6,
32'h03a90286,
32'h0296fe8b,
32'h011003dc,
32'h03780419,
32'h038e019a,
32'hfba30046,
32'hfc10fec0,
32'h015a027b,
32'h013fff87,
32'h026a0477,
32'hfe6803c0,
32'hfee9ff9e,
32'hfcfa020e,
32'hfc870320,
32'hfa37ff4e,
32'h0145fa7c,
32'h0351ff0c,
32'h01b40057,
32'hff1b0004,
32'hfc47022d,
32'hfde2fb80,
32'hfbe6fa8b,
32'hfc8e01bb,
32'hfe2a02f7,
32'h04d2fe9d,
32'h09540129,
32'h038f0366,
32'h03a9fbfd,
32'h0049ff77,
32'h013202de,
32'h0543ff15,
32'h00ff02a3,
32'h028302e7,
32'h005103a1,
32'h028102db,
32'h0546feb8,
32'h0115021f,
32'h0302053d,
32'hfcc90019,
32'hfe21f872,
32'h00b200d5,
32'hfa110679,
32'h00e6fb7f,
32'hfd44faf3,
32'hf807fbef,
32'h006cfd66,
32'h052701cc,
32'h068efd3b,
32'hff06fb2c,
32'hfd79fe9e,
32'h0365058a,
32'h01510359,
32'hfdfd0203,
32'h00fc04f9,
32'h093df71c,
32'h05c0fce1,
32'h000b07ae,
32'hfe9efd98,
32'hfbdf01f9,
32'h0165011c,
32'hffe5fd1e,
32'hffb501e5,
32'h019dfeee,
32'hfb4101a6,
32'hfef60265,
32'hfe040079,
32'hfa3e00f5,
32'hfa6ffdb2,
32'hfa5afb4b,
32'h0085f9da,
32'hfeaa006e,
32'h02500115,
32'h049efd57,
32'hfb3404cd,
32'hfe6803c0,
32'hfee9ff9e,
32'hfcfa020e,
32'hfc870320,
32'hfa37ff4e,
32'h0145fa7c,
32'h0351ff0c,
32'h01b40057,
32'hff1b0004,
32'hfc47022d,
32'hfde2fb80,
32'hfbe6fa8b,
32'hfc8e01bb,
32'hfe2a02f7,
32'h04d2fe9d,
32'h09540129,
32'h02e107ee,
32'hfedef96c,
32'h0294f4f0,
32'h01fb03e4,
32'h0044004d,
32'h0258fcf7,
32'h03f2003b,
32'h02160143,
32'hfe3a008c,
32'h01410305,
32'h001202ec,
32'hf4b8fd3c,
32'hf48f0078,
32'hfdcffc3d,
32'hfd81faa2,
32'hfd230558,
32'h051efddf,
32'h04defadd,
32'hffc70517,
32'h00ba00e0,
32'hfdb2fca5,
32'hfb5e0263,
32'hfed301c0,
32'h00940056,
32'h053d0540,
32'h06470072,
32'hff91fb0b,
32'hffacfae8,
32'hfe68fafb,
32'hf97502e3,
32'hfd05ffb1,
32'hfdf9fa40,
32'h00800080,
32'h047f0097,
32'hfdba00c5,
32'h01ad0120,
32'h0842000e,
32'h0138fb8a,
32'h0021fbdd,
32'h0196071c,
32'h03440223,
32'h0344ff4f,
32'hfc59013f,
32'hfd6bfa7c,
32'hffdb00de,
32'hfe70021f,
32'hfe33033a,
32'hfcc706e9,
32'hfe0002f0,
32'hfe8d08da,
32'h0094007e,
32'hff9ef78a,
32'hfb46fffe,
32'h01b001a3,
32'h02660561,
32'hfbe6031a,
32'hfe42fa8e,
32'h0185fb82,
32'h01d601bc,
32'hffe60349,
32'h01acfeef,
32'h040a032d,
32'h01f8fef4,
32'h04bdfd50,
32'h02e107ee,
32'hfedef96c,
32'h0294f4f0,
32'h01fb03e4,
32'h0044004d,
32'h0258fcf7,
32'h03f2003b,
32'h02160143,
32'hfe3a008c,
32'h01410305,
32'h001202ec,
32'hf4b8fd3c,
32'hf48f0078,
32'hfdcffc3d,
32'hfd81faa2,
32'hfd230558,
32'hff5ffa30,
32'h052d05aa,
32'h002005cf,
32'hfd990025,
32'hfddf0201,
32'hfe7e0508,
32'hfe61fde7,
32'hffa7f769,
32'hfd9efe18,
32'h00470042,
32'h04b7ff4e,
32'h03bafe2c,
32'h0654f73c,
32'hff45fd47,
32'hfc1e057a,
32'h0286ffcf,
32'hfd170259,
32'hfe540745,
32'h00e202ca,
32'hffda03c7,
32'h02f8031c,
32'hfa63fdbe,
32'hfa0bfed0,
32'h0311fdf5,
32'hffe2fd3e,
32'hfe58008f,
32'hff0cfd81,
32'hfc94fb3c,
32'hff29ffa3,
32'h01d90158,
32'hff01ff97,
32'h010fffc4,
32'h0390ffbf,
32'hff46fd4f,
32'h0043ff78,
32'hfee702bc,
32'hfacbffc3,
32'hfebcffff,
32'h038d02b3,
32'h06f10387,
32'h01320837,
32'hfab706f9,
32'hff88fef7,
32'h0034fd78,
32'hfee7fd78,
32'h00e6fd8c,
32'h01b4fe53,
32'h03feff54,
32'h06580476,
32'h03fffc22,
32'h00a8f481,
32'h02f50421,
32'h001e077e,
32'hfdb20057,
32'h03800050,
32'h0114fd0c,
32'hfe6c0171,
32'h0071fa6a,
32'h03c2f3e4,
32'h053f081e,
32'hfc590308,
32'hfb19f79f,
32'hfab2071f,
32'hf59801d8,
32'hff5ffa30,
32'h052d05aa,
32'h002005cf,
32'hfd990025,
32'hfddf0201,
32'hfe7e0508,
32'hfe61fde7,
32'hffa7f769,
32'hfd9efe18,
32'h00470042,
32'h04b7ff4e,
32'h03bafe2c,
32'h0654f73c,
32'hff45fd47,
32'hfc1e057a,
32'h0286ffcf,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f,
32'h0000000f};
