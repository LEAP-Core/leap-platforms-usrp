typedef        2048 NumSamples;
typedef        1363 PacketLength;

Bit#(32) samples[       2048] = {
32'hdeaddead,
32'hcafecafe,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h02f102f1,
32'h0026f786,
32'hfaf9ff23,
32'hff300922,
32'h000005e3,
32'hff300922,
32'hfaf9ff23,
32'h0026f786,
32'h02f102f1,
32'hf7860026,
32'hff23faf9,
32'h0922ff30,
32'h05e30000,
32'h0922ff30,
32'hff23faf9,
32'hf7860026,
32'h0000f600,
32'hf9c000c9,
32'hf93905de,
32'hf8a1fa1e,
32'hfc8fffd1,
32'h04bd04cd,
32'h014ff7d9,
32'h010ff832,
32'h09a8fdc1,
32'h0165fc62,
32'hfaccfc23,
32'hff180473,
32'hfa160543,
32'hfbd3f799,
32'hfd7cfc56,
32'hf9b4025c,
32'h04000400,
32'h004307a1,
32'hf5b7fe8f,
32'h00f403c1,
32'h03be0191,
32'h0308f73e,
32'h075c0010,
32'hffbd0369,
32'h01a8063e,
32'h06cbfd8c,
32'h0388f8a1,
32'h059d03d4,
32'hfe370159,
32'hfab30632,
32'h071d028b,
32'h07b3ffac,
32'h00000a00,
32'hf84cffac,
32'hf8e2028b,
32'h054c0632,
32'h01c80159,
32'hfa6203d4,
32'hfc77f8a1,
32'hf934fd8c,
32'hfe57063e,
32'h00420369,
32'hf8a30010,
32'hfcf7f73e,
32'hfc410191,
32'hff0b03c1,
32'h0a48fe8f,
32'hffbc07a1,
32'hfc000400,
32'h064b025c,
32'h0283fc56,
32'h042cf799,
32'h05e90543,
32'h00e70473,
32'h0533fc23,
32'hfe9afc62,
32'hf657fdc1,
32'hfef0f832,
32'hfeb0f7d9,
32'hfb4204cd,
32'h0370ffd1,
32'h075efa1e,
32'h06c605de,
32'h063f00c9,
32'h0000f600,
32'hf9c000c9,
32'hf93905de,
32'hf8a1fa1e,
32'hfc8fffd1,
32'h04bd04cd,
32'h014ff7d9,
32'h010ff832,
32'h09a8fdc1,
32'h0165fc62,
32'hfaccfc23,
32'hff180473,
32'hfa160543,
32'hfbd3f799,
32'hfd7cfc56,
32'hf9b4025c,
32'h04000400,
32'h004307a1,
32'hf5b7fe8f,
32'h00f403c1,
32'h03be0191,
32'h0308f73e,
32'h075c0010,
32'hffbd0369,
32'h01a8063e,
32'h06cbfd8c,
32'h0388f8a1,
32'h059d03d4,
32'hfe370159,
32'hfab30632,
32'h071d028b,
32'h07b3ffac,
32'h00000a00,
32'hf84cffac,
32'hf8e2028b,
32'h054c0632,
32'h01c80159,
32'hfa6203d4,
32'hfc77f8a1,
32'hf934fd8c,
32'hfe57063e,
32'h00420369,
32'hf8a30010,
32'hfcf7f73e,
32'hfc410191,
32'hff0b03c1,
32'h0a48fe8f,
32'hffbc07a1,
32'hfc000400,
32'h064b025c,
32'h0283fc56,
32'h042cf799,
32'h05e90543,
32'h00e70473,
32'h0533fc23,
32'hfe9afc62,
32'hf657fdc1,
32'hfef0f832,
32'hfeb0f7d9,
32'hfb4204cd,
32'h0370ffd1,
32'h075efa1e,
32'h06c605de,
32'h063f00c9,
32'h0000f600,
32'hf9c000c9,
32'hf93905de,
32'hf8a1fa1e,
32'hfc8fffd1,
32'h04bd04cd,
32'h014ff7d9,
32'h010ff832,
32'h09a8fdc1,
32'h0165fc62,
32'hfaccfc23,
32'hff180473,
32'hfa160543,
32'hfbd3f799,
32'hfd7cfc56,
32'hf9b4025c,
32'h04000400,
32'h004307a1,
32'hf5b7fe8f,
32'h00f403c1,
32'h03be0191,
32'h0308f73e,
32'h075c0010,
32'hffbd0369,
32'h01a8063e,
32'h06cbfd8c,
32'h0388f8a1,
32'h059d03d4,
32'hfe370159,
32'hfab30632,
32'h071d028b,
32'h07b3ffac,
32'hffff0200,
32'hfdfd083d,
32'hf84902f3,
32'hff8403c0,
32'h04f201e6,
32'h082cf89c,
32'h05bdfcf1,
32'hff01012c,
32'h03a7063d,
32'h01c8fc43,
32'h017ef9a2,
32'h088806a0,
32'hfbb7028d,
32'hfc43071c,
32'h0c960280,
32'h058bfdf5,
32'hfffd07fe,
32'hfa75fdf4,
32'hf36a027d,
32'h03bb071c,
32'h0446028d,
32'hf775069d,
32'hfe81f9a1,
32'hfe39fc45,
32'hfc57063d,
32'h00fd012c,
32'hfa40fcf0,
32'hf7d4f898,
32'hfb0e01e6,
32'h007a03c0,
32'h07b602f4,
32'h0200083e,
32'h000001ff,
32'h053c03f8,
32'h03a5f97b,
32'h04d5f3ad,
32'h01e107c2,
32'hffaf03e0,
32'h0549fb90,
32'hfd1b01f3,
32'hf858fdc0,
32'h01bcf627,
32'hff32fa8c,
32'hfc42013a,
32'h031bfbca,
32'h0506fd21,
32'h04ff0462,
32'h05140047,
32'h0000fc00,
32'hfaeb0047,
32'hfaff0461,
32'hfafbfd21,
32'hfce4fbcb,
32'h03bc0139,
32'h00cefa8d,
32'hfe44f626,
32'h07a7fdc3,
32'h02e401f6,
32'hfab6fb8f,
32'h005003e0,
32'hfe1e07c1,
32'hfb2ef3ac,
32'hfc5bf97b,
32'hfac303f8,
32'hffff0200,
32'hfdfd083d,
32'hf84902f3,
32'hff8403c0,
32'h04f201e6,
32'h082cf89c,
32'h05bdfcf1,
32'hff01012c,
32'h03a7063d,
32'h01c8fc43,
32'h017ef9a2,
32'h088806a0,
32'hfbb7028d,
32'hfc43071c,
32'h0c960280,
32'h058bfdf5,
32'hfb5f011e,
32'hf951017d,
32'h019000c7,
32'hfddcfeea,
32'hfb790386,
32'hfa39037b,
32'hf786fe70,
32'hfdaefe19,
32'h0008fc85,
32'hf936fd36,
32'hfba6ffa0,
32'h065b0130,
32'h011c0477,
32'hfa3d019f,
32'hffb000fe,
32'hfe760296,
32'hfdc9fd76,
32'h012af98f,
32'h0194faf6,
32'h02580463,
32'h008d0370,
32'hfeb6f768,
32'hff2efe0f,
32'h023b06e9,
32'h017b01de,
32'hfe3bfbcf,
32'hff36facc,
32'hfd2a0002,
32'h02740112,
32'h0620ffd9,
32'hfcdb0239,
32'hff790130,
32'h0290fe50,
32'hfe3efd59,
32'h0478fd92,
32'h060afe38,
32'hfbc802e5,
32'hfd2c0668,
32'h05800491,
32'hfd340358,
32'hfdc8ff0a,
32'h08ddffb8,
32'h010c0387,
32'h0322fe1c,
32'h0729fc49,
32'hf900fe38,
32'hfc87006b,
32'h070502e1,
32'h03c60378,
32'hff7c0583,
32'hfdc2fdb1,
32'hffd5f7a2,
32'h014ffb61,
32'hff30f9f0,
32'h0046ff9a,
32'h053905b9,
32'h033300f1,
32'hfd6dfebe,
32'hfdf7fe89,
32'h00d70183,
32'h05a402af,
32'h0362fdaa,
32'hffb0ffae,
32'h031b034a,
32'hfb5f011e,
32'hf951017d,
32'h019000c7,
32'hfddcfeea,
32'hfb790386,
32'hfa39037b,
32'hf786fe70,
32'hfdaefe19,
32'h0008fc85,
32'hf936fd36,
32'hfba6ffa0,
32'h065b0130,
32'h011c0477,
32'hfa3d019f,
32'hffb000fe,
32'hfe760296,
32'h004605c7,
32'h040bfe1c,
32'hfebffe4b,
32'hfda9fbca,
32'hfed100a8,
32'hfdda05f4,
32'hfca7ff7d,
32'h0495027d,
32'h06460012,
32'hf8defbbd,
32'hfe77062f,
32'h0690051f,
32'hff3b001b,
32'h02d7035c,
32'h0444006f,
32'hfac4fae0,
32'hfba1f8de,
32'h02e40191,
32'h02b706e6,
32'h009c003f,
32'hff640378,
32'hfdb10177,
32'hffc1fbda,
32'h0195034b,
32'h04c200fe,
32'h039d0093,
32'h004102b6,
32'h0618fc82,
32'h015902f8,
32'hfd6e0512,
32'h0192025c,
32'hfbf9040d,
32'h00d8fc17,
32'h0208fbb4,
32'hfdf3fc63,
32'h060cf8e4,
32'hfd0ffd13,
32'hf74cfbcb,
32'h025afe19,
32'h01c2045b,
32'hff2803bd,
32'hff3800da,
32'hfe93fd66,
32'hffbd0032,
32'hff9bfe21,
32'hfd1bfc59,
32'hfcda0651,
32'h0407049a,
32'h04bf00c0,
32'hff8205fd,
32'hfe540396,
32'hfaa4fe9a,
32'hfafcfc4a,
32'hfe70f9ca,
32'hfc1bfad8,
32'hfdf1ff9e,
32'h01cdff72,
32'hfaeffda2,
32'hfc34fe86,
32'h08f4fc13,
32'h030f018b,
32'hfdb70285,
32'h0432f89a,
32'hff8900ca,
32'h004605c7,
32'h040bfe1c,
32'hfebffe4b,
32'hfda9fbca,
32'hfed100a8,
32'hfdda05f4,
32'hfca7ff7d,
32'h0495027d,
32'h06460012,
32'hf8defbbd,
32'hfe77062f,
32'h0690051f,
32'hff3b001b,
32'h02d7035c,
32'h0444006f,
32'hfac4fae0,
32'hfd50feb7,
32'h00fdfdfd,
32'h0668004f,
32'hfec0063a,
32'hfcf6064b,
32'h0112fc86,
32'hfbaef7ea,
32'h01a3fd27,
32'h03360329,
32'hfea30320,
32'h012900ce,
32'h002d00d1,
32'h0374009f,
32'h02e5fed5,
32'hfdb2fe1d,
32'hfcfafefa,
32'hff00ff36,
32'h011dfc82,
32'hfad7f97c,
32'hfd340083,
32'h007e0446,
32'hfafbff14,
32'hfe640844,
32'hfae7089d,
32'hfa6ff67f,
32'h020ff531,
32'h0014fe81,
32'h01ee0672,
32'h031907c2,
32'h0096ff84,
32'hfd71fcb5,
32'h0000fdf8,
32'h089f00d9,
32'hfe28033d,
32'hf9430088,
32'h01affc65,
32'hfa08fcfa,
32'hf95f02bb,
32'h019cfec1,
32'hffc9fc86,
32'hfef800c7,
32'h0247fd99,
32'h042a02eb,
32'h051a01c1,
32'h0697f988,
32'h0418035f,
32'h01ca0627,
32'h05080133,
32'h01af01b7,
32'hfc5300b3,
32'h03c30118,
32'h05f0fde4,
32'hfc82fbd1,
32'h002bfe1c,
32'h031afea6,
32'hfbd7fe68,
32'hfec3004f,
32'hfff70557,
32'hff1001da,
32'hff93ff6d,
32'hfc5904f5,
32'h014b001e,
32'h0207fc6e,
32'hfd6fffab,
32'hfd50feb7,
32'h00fdfdfd,
32'h0668004f,
32'hfec0063a,
32'hfcf6064b,
32'h0112fc86,
32'hfbaef7ea,
32'h01a3fd27,
32'h03360329,
32'hfea30320,
32'h012900ce,
32'h002d00d1,
32'h0374009f,
32'h02e5fed5,
32'hfdb2fe1d,
32'hfcfafefa,
32'h064f0268,
32'h02000196,
32'h03c3ff76,
32'hfef7fc1d,
32'hfbe3ffba,
32'hff92ff02,
32'h00980257,
32'hfffd02bb,
32'hfc07fc24,
32'h01adfd13,
32'h01660132,
32'hfced029a,
32'h01d7fdae,
32'hffe1ff7f,
32'h015306ff,
32'h01b805e3,
32'h003f04c6,
32'h02d1ff28,
32'hff76fd81,
32'h004c00bf,
32'hfe9cfac6,
32'hff90fd29,
32'h0266ff08,
32'hfedffe61,
32'h05f30670,
32'h01270086,
32'hf9eefbe4,
32'h048b0555,
32'h022603ca,
32'hfa23fd8e,
32'hfab5fdce,
32'hffb1ff44,
32'h03d00058,
32'h01a6fd9d,
32'hfe41fd3c,
32'hfbc80412,
32'h017202de,
32'h0374fc6e,
32'hfd5dfe2f,
32'h0047ff18,
32'h0209fecb,
32'h01b3015d,
32'h07d40205,
32'h06e5008f,
32'hfb92feb8,
32'hfce3ff4d,
32'h0670fe96,
32'h0369fd89,
32'h03a0fcf8,
32'hfee3fbe1,
32'hf75b005f,
32'h0037ffe0,
32'hfecefd20,
32'hf9fb0234,
32'hfbbc0513,
32'hfbfe0305,
32'hff3cf99f,
32'hfdc6f6ee,
32'h00ff000f,
32'hfe3d0198,
32'hf9ef004d,
32'h02ddffb3,
32'hfeec03b7,
32'h0027082c,
32'h064f0268,
32'h02000196,
32'h03c3ff76,
32'hfef7fc1d,
32'hfbe3ffba,
32'hff92ff02,
32'h00980257,
32'hfffd02bb,
32'hfc07fc24,
32'h01adfd13,
32'h01660132,
32'hfced029a,
32'h01d7fdae,
32'hffe1ff7f,
32'h015306ff,
32'h01b805e3,
32'h010f0380,
32'hfcb20009,
32'h026bfa37,
32'h028efd50,
32'hfc36feab,
32'hffd6fa98,
32'h0152fcee,
32'h0001048f,
32'h01a20714,
32'hff84ff6d,
32'hfffaf9b2,
32'h05e4fc3d,
32'h058afa34,
32'hfe1ffd12,
32'hfb6e0252,
32'hfcc5fccf,
32'hfc080086,
32'hfd8a02c2,
32'h00dbfd50,
32'h01840083,
32'h0295fc7a,
32'h06c4f97a,
32'h0694fdb9,
32'h015afe64,
32'h00f501d8,
32'h00d20212,
32'h00da0030,
32'h053ffcdc,
32'h021afb59,
32'hfa28ff59,
32'hf8ef0055,
32'hfb2e04ce,
32'hfbbf034f,
32'hfd100727,
32'h00441149,
32'hff16004e,
32'hfddffaf3,
32'hfe6a055d,
32'hfda5fffc,
32'h03530156,
32'h02bdfdab,
32'hfa94f971,
32'h012901a2,
32'h05470166,
32'hfc610083,
32'hffa8fdf3,
32'h059afadf,
32'hfcba01b0,
32'hfca60727,
32'h063c0416,
32'h016afefc,
32'hff0f034f,
32'h061504a6,
32'h01b30247,
32'hfda606d4,
32'hfece02f8,
32'hf9aa00a6,
32'hfb7c0005,
32'h018cf76d,
32'hfe5ffd2a,
32'hffba04ef,
32'h0367fe68,
32'hff53fac0,
32'h00cdfed3,
32'h010f0380,
32'hfcb20009,
32'h026bfa37,
32'h028efd50,
32'hfc36feab,
32'hffd6fa98,
32'h0152fcee,
32'h0001048f,
32'h01a20714,
32'hff84ff6d,
32'hfffaf9b2,
32'h05e4fc3d,
32'h058afa34,
32'hfe1ffd12,
32'hfb6e0252,
32'hfcc5fccf,
32'h0320fc21,
32'h043101a0,
32'h00b50019,
32'hf730fd52,
32'hfa15fede,
32'hfd7afbd2,
32'h00befafa,
32'h007402e5,
32'hfc37051f,
32'h032cfe56,
32'h012a0156,
32'hfd760821,
32'h05c2038c,
32'h07170041,
32'h0186024c,
32'hfdb0060a,
32'hfb460695,
32'hf9c3014f,
32'h01db00c6,
32'h0166fb29,
32'hf877f70d,
32'h028102db,
32'h00cf0471,
32'hfc0d005a,
32'h05fe03bf,
32'hffd9ff8b,
32'hfeaafec0,
32'hffa5025a,
32'hf9b5ff86,
32'h003d0028,
32'h01cdfd1c,
32'hffaaf6ec,
32'hffe0fe40,
32'h039503db,
32'h073402d8,
32'hfe7d0663,
32'h002303e4,
32'h061aff80,
32'h009ffaf4,
32'h00c8f83b,
32'h009704cf,
32'hfd6504d3,
32'h014cf7c4,
32'h02effa80,
32'hff2a00ea,
32'h036d063d,
32'h031b01fc,
32'hf913f897,
32'hfe38fe87,
32'h02fbfeb7,
32'hfebafcea,
32'h023b025b,
32'h0231fd4d,
32'hfd16fcc0,
32'hfd3102df,
32'h046100cd,
32'h05f2fa12,
32'hfe12f62b,
32'hfbdffe01,
32'hfeac04ee,
32'h043b0123,
32'h000a0384,
32'hf7b10758,
32'hfedcff80,
32'h0320fc21,
32'h043101a0,
32'h00b50019,
32'hf730fd52,
32'hfa15fede,
32'hfd7afbd2,
32'h00befafa,
32'h007402e5,
32'hfc37051f,
32'h032cfe56,
32'h012a0156,
32'hfd760821,
32'h05c2038c,
32'h07170041,
32'h0186024c,
32'hfdb0060a,
32'h010606a0,
32'h061803ba,
32'h01abf970,
32'hfc340065,
32'h0116febd,
32'h038cfdf6,
32'h00bd0347,
32'hfdfcfb89,
32'h02f4ffba,
32'h00c300eb,
32'hfa21ff67,
32'hffd5048f,
32'h00ca0234,
32'h03e9076d,
32'h082b025f,
32'hff1afed5,
32'hfb47055d,
32'hfebafc29,
32'h021fff8a,
32'hffbd0235,
32'hfab3fd07,
32'hfbc40323,
32'hfd98fe18,
32'h017afc03,
32'hff42fe4c,
32'hfda2fc80,
32'hfd99009f,
32'hf3b7fd7e,
32'hfb96ffe5,
32'h04530954,
32'hfca704ad,
32'h0054ffe0,
32'h03080290,
32'h01dcfd1c,
32'hff97f768,
32'hfa8ffce2,
32'hff40fe5e,
32'h02d5ff0f,
32'h030f02e3,
32'hfeb10226,
32'hfb5b0315,
32'h029f0173,
32'hff35001c,
32'hfa8dff86,
32'h010ffdd8,
32'h0206009d,
32'h0254ff9f,
32'h032b02ba,
32'hfe67038f,
32'hfddbff26,
32'h01a30456,
32'hff83ff65,
32'h0138f73c,
32'h0840fa86,
32'h0444fe0a,
32'h0288ff75,
32'h06aefc44,
32'hfecdfeb6,
32'hfa4a0261,
32'h02a6febb,
32'h014ffdae,
32'hf9f5ffb7,
32'hffec0148,
32'h02f100b2,
32'h010606a0,
32'h061803ba,
32'h01abf970,
32'hfc340065,
32'h0116febd,
32'h038cfdf6,
32'h00bd0347,
32'hfdfcfb89,
32'h02f4ffba,
32'h00c300eb,
32'hfa21ff67,
32'hffd5048f,
32'h00ca0234,
32'h03e9076d,
32'h082b025f,
32'hff1afed5,
32'h0358fc90,
32'hf977fca6,
32'hfbfefe1e,
32'h0c2bfbf1,
32'h02a6fc33,
32'hfb04ffe2,
32'h0021015b,
32'hfe0a0506,
32'hfd20064c,
32'h029ffe3f,
32'h0782fb6c,
32'hffb0ff7f,
32'hfbbffd80,
32'hfe3dfb30,
32'hfc76fdc4,
32'h016bfcc0,
32'hfc60fe36,
32'hf9b10540,
32'h0340035b,
32'h0265ffec,
32'h027900ac,
32'hfd69fd6b,
32'hfd43fea4,
32'h085b0030,
32'h040dff88,
32'h014c068a,
32'h003c04a7,
32'hfd4df813,
32'h00d8f8c0,
32'hff4e0116,
32'h002b024a,
32'hff6a0104,
32'h021701d0,
32'h06000572,
32'hfb280403,
32'hfe4cfd49,
32'h05cfff47,
32'hfbb0fef1,
32'hf7b0fc09,
32'hfe3d02dd,
32'h01ae0192,
32'hf94afdb4,
32'hfa6100cb,
32'h0757ff94,
32'h00b2fd32,
32'hfcaafbbd,
32'h04cf010e,
32'h00cf00bf,
32'h0231f928,
32'h06160174,
32'hfd4400f2,
32'hfdbffcab,
32'hffce0899,
32'hfb18062c,
32'h0368026f,
32'h07730607,
32'hfee10157,
32'hfac600fb,
32'hfb33fd6e,
32'h0198fa5c,
32'h0636024c,
32'h02d504c4,
32'hfd0f02a8,
32'hfe38008b,
32'h0358fc90,
32'hf977fca6,
32'hfbfefe1e,
32'h0c2bfbf1,
32'h02a6fc33,
32'hfb04ffe2,
32'h0021015b,
32'hfe0a0506,
32'hfd20064c,
32'h029ffe3f,
32'h0782fb6c,
32'hffb0ff7f,
32'hfbbffd80,
32'hfe3dfb30,
32'hfc76fdc4,
32'h016bfcc0,
32'h05df00b9,
32'h00dfffa2,
32'hffcff85d,
32'h0752fed3,
32'hfcec000d,
32'hfcf6fff7,
32'h028603a9,
32'hfe8b0296,
32'h03dc0110,
32'h04190378,
32'h019a038e,
32'h0046fba3,
32'hfec0fc10,
32'h027b015a,
32'hff87013f,
32'h0477026a,
32'h028fff07,
32'hf6dd015b,
32'h007e02f8,
32'hffadfaba,
32'hf9e0fb03,
32'hfee7f807,
32'hfd8ef888,
32'h04d70599,
32'h05d6049a,
32'h005cfe65,
32'h016b0072,
32'h00b600bb,
32'h050000ad,
32'h01c2006e,
32'h012ffcdf,
32'h04670102,
32'hfbde0806,
32'h0140051e,
32'h03e3046b,
32'hfb70ffdb,
32'h0055fc82,
32'h011b0669,
32'hfe34010b,
32'h014ff891,
32'hff43fbf0,
32'hfe86fcc1,
32'h01850154,
32'hf7a500f1,
32'hf2140089,
32'h00690214,
32'hfe58fe4e,
32'hf6e603c8,
32'hfed00237,
32'hfb38fc17,
32'hfc1700cc,
32'h02a3fe8f,
32'hff7ffc6c,
32'h02490311,
32'h019f061b,
32'h01340063,
32'h02a8fe26,
32'hfca20301,
32'h0329ff1c,
32'h048cfb37,
32'hf9cb0276,
32'h013e0752,
32'h0407fdba,
32'hff0ff6a6,
32'h05df00b9,
32'h00dfffa2,
32'hffcff85d,
32'h0752fed3,
32'hfcec000d,
32'hfcf6fff7,
32'h028603a9,
32'hfe8b0296,
32'h03dc0110,
32'h04190378,
32'h019a038e,
32'h0046fba3,
32'hfec0fc10,
32'h027b015a,
32'hff87013f,
32'h0477026a,
32'h03c0fe68,
32'hff9efee9,
32'h020efcfa,
32'h0320fc87,
32'hff4efa37,
32'hfa7c0145,
32'hff0c0351,
32'h005701b4,
32'h0004ff1b,
32'h022dfc47,
32'hfb80fde2,
32'hfa8bfbe6,
32'h01bbfc8e,
32'h02f7fe2a,
32'hfe9d04d2,
32'h01290954,
32'h0366038f,
32'hfbfd03a9,
32'hff770049,
32'h02de0132,
32'hff150543,
32'h02a300ff,
32'h02e70283,
32'h03a10051,
32'h02db0281,
32'hfeb80546,
32'h021f0115,
32'h053d0302,
32'h0019fcc9,
32'hf872fe21,
32'h00d500b2,
32'h0679fa11,
32'hfb7f00e6,
32'hfaf3fd44,
32'hfbeff807,
32'hfd66006c,
32'h01cc0527,
32'hfd3b068e,
32'hfb2cff06,
32'hfe9efd79,
32'h058a0365,
32'h03590151,
32'h0203fdfd,
32'h04f900fc,
32'hf71c093d,
32'hfce105c0,
32'h07ae000b,
32'hfd98fe9e,
32'h01f9fbdf,
32'h011c0165,
32'hfd1effe5,
32'h01e5ffb5,
32'hfeee019d,
32'h01a6fb41,
32'h0265fef6,
32'h0079fe04,
32'h00f5fa3e,
32'hfdb2fa6f,
32'hfb4bfa5a,
32'hf9da0085,
32'h006efeaa,
32'h01150250,
32'hfd57049e,
32'h04cdfb34,
32'h03c0fe68,
32'hff9efee9,
32'h020efcfa,
32'h0320fc87,
32'hff4efa37,
32'hfa7c0145,
32'hff0c0351,
32'h005701b4,
32'h0004ff1b,
32'h022dfc47,
32'hfb80fde2,
32'hfa8bfbe6,
32'h01bbfc8e,
32'h02f7fe2a,
32'hfe9d04d2,
32'h01290954,
32'h07ee02e1,
32'hf96cfede,
32'hf4f00294,
32'h03e401fb,
32'h004d0044,
32'hfcf70258,
32'h003b03f2,
32'h01430216,
32'h008cfe3a,
32'h03050141,
32'h02ec0012,
32'hfd3cf4b8,
32'h0078f48f,
32'hfc3dfdcf,
32'hfaa2fd81,
32'h0558fd23,
32'hfddf051e,
32'hfadd04de,
32'h0517ffc7,
32'h00e000ba,
32'hfca5fdb2,
32'h0263fb5e,
32'h01c0fed3,
32'h00560094,
32'h0540053d,
32'h00720647,
32'hfb0bff91,
32'hfae8ffac,
32'hfafbfe68,
32'h02e3f975,
32'hffb1fd05,
32'hfa40fdf9,
32'h00800080,
32'h0097047f,
32'h00c5fdba,
32'h012001ad,
32'h000e0842,
32'hfb8a0138,
32'hfbdd0021,
32'h071c0196,
32'h02230344,
32'hff4f0344,
32'h013ffc59,
32'hfa7cfd6b,
32'h00deffdb,
32'h021ffe70,
32'h033afe33,
32'h06e9fcc7,
32'h02f0fe00,
32'h08dafe8d,
32'h007e0094,
32'hf78aff9e,
32'hfffefb46,
32'h01a301b0,
32'h05610266,
32'h031afbe6,
32'hfa8efe42,
32'hfb820185,
32'h01bc01d6,
32'h0349ffe6,
32'hfeef01ac,
32'h032d040a,
32'hfef401f8,
32'hfd5004bd,
32'h07ee02e1,
32'hf96cfede,
32'hf4f00294,
32'h03e401fb,
32'h004d0044,
32'hfcf70258,
32'h003b03f2,
32'h01430216,
32'h008cfe3a,
32'h03050141,
32'h02ec0012,
32'hfd3cf4b8,
32'h0078f48f,
32'hfc3dfdcf,
32'hfaa2fd81,
32'h0558fd23,
32'hfa30ff5f,
32'h05aa052d,
32'h05cf0020,
32'h0025fd99,
32'h0201fddf,
32'h0508fe7e,
32'hfde7fe61,
32'hf769ffa7,
32'hfe18fd9e,
32'h00420047,
32'hff4e04b7,
32'hfe2c03ba,
32'hf73c0654,
32'hfd47ff45,
32'h057afc1e,
32'hffcf0286,
32'h0259fd17,
32'h0745fe54,
32'h02ca00e2,
32'h03c7ffda,
32'h031c02f8,
32'hfdbefa63,
32'hfed0fa0b,
32'hfdf50311,
32'hfd3effe2,
32'h008ffe58,
32'hfd81ff0c,
32'hfb3cfc94,
32'hffa3ff29,
32'h015801d9,
32'hff97ff01,
32'hffc4010f,
32'hffbf0390,
32'hfd4fff46,
32'hff780043,
32'h02bcfee7,
32'hffc3facb,
32'hfffffebc,
32'h02b3038d,
32'h038706f1,
32'h08370132,
32'h06f9fab7,
32'hfef7ff88,
32'hfd780034,
32'hfd78fee7,
32'hfd8c00e6,
32'hfe5301b4,
32'hff5403fe,
32'h04760658,
32'hfc2203ff,
32'hf48100a8,
32'h042102f5,
32'h077e001e,
32'h0057fdb2,
32'h00500380,
32'hfd0c0114,
32'h0171fe6c,
32'hfa6a0071,
32'hf3e403c2,
32'h081e053f,
32'h0308fc59,
32'hf79ffb19,
32'h071ffab2,
32'h01d8f598,
32'hfa30ff5f,
32'h05aa052d,
32'h05cf0020,
32'h0025fd99,
32'h0201fddf,
32'h0508fe7e,
32'hfde7fe61,
32'hf769ffa7,
32'hfe18fd9e,
32'h00420047,
32'hff4e04b7,
32'hfe2c03ba,
32'hf73c0654,
32'hfd47ff45,
32'h057afc1e,
32'hffcf0286,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h000f0000,
32'h0000000f};
